CDLv2�H�\                                                                                                                   		                             		  		                                                                                                     	          	                                                                                                                                                                                                                                                                                                        	                                    	                                                             	                                    		        	          				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                							      				                      	   	                                                                                                   	                                 				                                                                                                                                                             	   		                                                                       	                                                                                                                                                                          			                                                                                                                                                                                                                                                       	                                          						             				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              			                                                                                                                                  	     				                         	                                       	                                     			                    	                                                                                      	                     	                                                                                                                                                     	                                                                                                                                                                                                                                                                     	                                                                                                                                                                                                                                                                                                                                                                             	  	                     		          			                       			             						                                        	                                                                              	                                                                                                                                                                                                                   	                                                                                                                                         	                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                               		    	                                                                	                                                                               	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	            	            	                                                        	                                                                                      	            	                                                                      		       		          		                                                                       	                                                    					                                    	                              		                   	 	       	 			   	      	                                               			                                           	                        			                    			      		   		                  	                     				                                                                                                                            	                                                                                                                                         					    	          	                                                                                                                                                                                                                              	                                                                                                                                                                                           					        			                                                                                                                                                                                                   	                                                			                  				          							          	 					 	      	                                                                                             									                                                 		                                                                	                        	                       			    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         